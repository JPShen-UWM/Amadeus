module weight_buffer(
    input clk,
    input rst_n,
    in
);


endmodule