module weight_buffer(
    input clk,
    input rst_n,
    input start,
    input op_mode,
    input mem_ack,
    input [63:0] weight_data,
    output mem_req
);


endmodule