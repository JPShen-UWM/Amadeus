module ifmp_buffer(
    input clk,
    input rst_n,
    

);


endmodule