`include "sv/sys_defs.svh"

class 