module psum_buffer(
    input clk,
    input rst_n,
    input start,
    input start_conv
    output 
);
    


endmodule