module ifmap_buffer(
    input clk,
    input rst_n,
    input DECOMRPESS_FIFO_PACKET decompressed_fifo_packet,
    output 
);

endmodule