// Processing element