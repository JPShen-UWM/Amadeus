module NOC(
    input clk,
    input rst_n,
    input start,
    input LAYER_TYPE layer_type_in,
    input 
    output 
    output free_ifmap_buffer
);
    
    

endmodule